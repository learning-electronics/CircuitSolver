*Simple linear example

example exercise
V1 1 0 2V
R1 1 2 2ohm
R2 2 3 2ohm
Vm 4 3 0
R3 4 5 2ohm
R4 5 6 2ohm
H1 6 0 Vm 2
.END
