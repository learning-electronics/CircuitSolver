*Simple linear example

example exercise
R1 1 0 1Kohm
V1 1 0 5V
V2 1 2 6V
C1 2 0 1UF
.END
