*Simple linear example

example exercise
V1 4 1 2V
V2 4 2 
.END
