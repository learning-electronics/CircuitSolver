*Simple linear example

example exercise
R1 2 1 4ohm
R2 1 0 2ohm
V1 2 0 6V
.END
